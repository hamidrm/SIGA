----------------------------------------------------------------------------------
-- SIGA
-- Author: Hamidreza Mehrabian
-- File: siga_utilities.vhdl
-- Description: a package for types and functions
----------------------------------------------------------------------------------
library IEEE;

use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
package siga_utilities is

-------------------------------------------------------------------------
-- Types
-------------------------------------------------------------------------

type mem_mul_r_14b_t is array (0 to 599) of std_logic_vector(13 downto 0);
type siga_re_cmd_t is (RASTER_FILL_RECT, RASTER_DRAW_LINE, RASTER_DRAW_CIRCLE, RASTER_FILL_CIRCLE, RASTER_FILL_RECT_BMP);
subtype siga_re_params_t is integer range -800 to 800;

type siga_point2_t is
record
x : std_logic_vector(9 downto 0); -- [0 to 799]
y : std_logic_vector(9 downto 0); -- [0 to 599]
end record;

type siga_rgb_t is
record
r : std_logic_vector(4 downto 0);
g : std_logic_vector(5 downto 0);
b : std_logic_vector(4 downto 0);
end record;

type siga_fb_cmd_t is
record
color       : siga_rgb_t;                   -- Color in RGB 5:6:5
fill_length : std_logic_vector(7 downto 0); -- Length of burst filling
pos         : siga_point2_t;                -- Coordinate of start point
dest_addr   : std_logic_vector(3 downto 0); -- Most significant 3 bits of the destination buffer address
--solid_color        		: std_logic; 							 -- Is this command a solid color?
end record;
-------------------------------------------------------------------------
-- Constants
-------------------------------------------------------------------------
constant mul_r_c_table : mem_mul_r_14b_t := (
	"00000000000000",
	"00000000011001",
	"00000000110010",
	"00000001001011",
	"00000001100100",
	"00000001111101",
	"00000010010110",
	"00000010101111",
	"00000011001000",
	"00000011100001",
	"00000011111010",
	"00000100010011",
	"00000100101100",
	"00000101000101",
	"00000101011110",
	"00000101110111",
	"00000110010000",
	"00000110101001",
	"00000111000010",
	"00000111011011",
	"00000111110100",
	"00001000001101",
	"00001000100110",
	"00001000111111",
	"00001001011000",
	"00001001110001",
	"00001010001010",
	"00001010100011",
	"00001010111100",
	"00001011010101",
	"00001011101110",
	"00001100000111",
	"00001100100000",
	"00001100111001",
	"00001101010010",
	"00001101101011",
	"00001110000100",
	"00001110011101",
	"00001110110110",
	"00001111001111",
	"00001111101000",
	"00010000000001",
	"00010000011010",
	"00010000110011",
	"00010001001100",
	"00010001100101",
	"00010001111110",
	"00010010010111",
	"00010010110000",
	"00010011001001",
	"00010011100010",
	"00010011111011",
	"00010100010100",
	"00010100101101",
	"00010101000110",
	"00010101011111",
	"00010101111000",
	"00010110010001",
	"00010110101010",
	"00010111000011",
	"00010111011100",
	"00010111110101",
	"00011000001110",
	"00011000100111",
	"00011001000000",
	"00011001011001",
	"00011001110010",
	"00011010001011",
	"00011010100100",
	"00011010111101",
	"00011011010110",
	"00011011101111",
	"00011100001000",
	"00011100100001",
	"00011100111010",
	"00011101010011",
	"00011101101100",
	"00011110000101",
	"00011110011110",
	"00011110110111",
	"00011111010000",
	"00011111101001",
	"00100000000010",
	"00100000011011",
	"00100000110100",
	"00100001001101",
	"00100001100110",
	"00100001111111",
	"00100010011000",
	"00100010110001",
	"00100011001010",
	"00100011100011",
	"00100011111100",
	"00100100010101",
	"00100100101110",
	"00100101000111",
	"00100101100000",
	"00100101111001",
	"00100110010010",
	"00100110101011",
	"00100111000100",
	"00100111011101",
	"00100111110110",
	"00101000001111",
	"00101000101000",
	"00101001000001",
	"00101001011010",
	"00101001110011",
	"00101010001100",
	"00101010100101",
	"00101010111110",
	"00101011010111",
	"00101011110000",
	"00101100001001",
	"00101100100010",
	"00101100111011",
	"00101101010100",
	"00101101101101",
	"00101110000110",
	"00101110011111",
	"00101110111000",
	"00101111010001",
	"00101111101010",
	"00110000000011",
	"00110000011100",
	"00110000110101",
	"00110001001110",
	"00110001100111",
	"00110010000000",
	"00110010011001",
	"00110010110010",
	"00110011001011",
	"00110011100100",
	"00110011111101",
	"00110100010110",
	"00110100101111",
	"00110101001000",
	"00110101100001",
	"00110101111010",
	"00110110010011",
	"00110110101100",
	"00110111000101",
	"00110111011110",
	"00110111110111",
	"00111000010000",
	"00111000101001",
	"00111001000010",
	"00111001011011",
	"00111001110100",
	"00111010001101",
	"00111010100110",
	"00111010111111",
	"00111011011000",
	"00111011110001",
	"00111100001010",
	"00111100100011",
	"00111100111100",
	"00111101010101",
	"00111101101110",
	"00111110000111",
	"00111110100000",
	"00111110111001",
	"00111111010010",
	"00111111101011",
	"01000000000100",
	"01000000011101",
	"01000000110110",
	"01000001001111",
	"01000001101000",
	"01000010000001",
	"01000010011010",
	"01000010110011",
	"01000011001100",
	"01000011100101",
	"01000011111110",
	"01000100010111",
	"01000100110000",
	"01000101001001",
	"01000101100010",
	"01000101111011",
	"01000110010100",
	"01000110101101",
	"01000111000110",
	"01000111011111",
	"01000111111000",
	"01001000010001",
	"01001000101010",
	"01001001000011",
	"01001001011100",
	"01001001110101",
	"01001010001110",
	"01001010100111",
	"01001011000000",
	"01001011011001",
	"01001011110010",
	"01001100001011",
	"01001100100100",
	"01001100111101",
	"01001101010110",
	"01001101101111",
	"01001110001000",
	"01001110100001",
	"01001110111010",
	"01001111010011",
	"01001111101100",
	"01010000000101",
	"01010000011110",
	"01010000110111",
	"01010001010000",
	"01010001101001",
	"01010010000010",
	"01010010011011",
	"01010010110100",
	"01010011001101",
	"01010011100110",
	"01010011111111",
	"01010100011000",
	"01010100110001",
	"01010101001010",
	"01010101100011",
	"01010101111100",
	"01010110010101",
	"01010110101110",
	"01010111000111",
	"01010111100000",
	"01010111111001",
	"01011000010010",
	"01011000101011",
	"01011001000100",
	"01011001011101",
	"01011001110110",
	"01011010001111",
	"01011010101000",
	"01011011000001",
	"01011011011010",
	"01011011110011",
	"01011100001100",
	"01011100100101",
	"01011100111110",
	"01011101010111",
	"01011101110000",
	"01011110001001",
	"01011110100010",
	"01011110111011",
	"01011111010100",
	"01011111101101",
	"01100000000110",
	"01100000011111",
	"01100000111000",
	"01100001010001",
	"01100001101010",
	"01100010000011",
	"01100010011100",
	"01100010110101",
	"01100011001110",
	"01100011100111",
	"01100100000000",
	"01100100011001",
	"01100100110010",
	"01100101001011",
	"01100101100100",
	"01100101111101",
	"01100110010110",
	"01100110101111",
	"01100111001000",
	"01100111100001",
	"01100111111010",
	"01101000010011",
	"01101000101100",
	"01101001000101",
	"01101001011110",
	"01101001110111",
	"01101010010000",
	"01101010101001",
	"01101011000010",
	"01101011011011",
	"01101011110100",
	"01101100001101",
	"01101100100110",
	"01101100111111",
	"01101101011000",
	"01101101110001",
	"01101110001010",
	"01101110100011",
	"01101110111100",
	"01101111010101",
	"01101111101110",
	"01110000000111",
	"01110000100000",
	"01110000111001",
	"01110001010010",
	"01110001101011",
	"01110010000100",
	"01110010011101",
	"01110010110110",
	"01110011001111",
	"01110011101000",
	"01110100000001",
	"01110100011010",
	"01110100110011",
	"01110101001100",
	"01110101100101",
	"01110101111110",
	"01110110010111",
	"01110110110000",
	"01110111001001",
	"01110111100010",
	"01110111111011",
	"01111000010100",
	"01111000101101",
	"01111001000110",
	"01111001011111",
	"01111001111000",
	"01111010010001",
	"01111010101010",
	"01111011000011",
	"01111011011100",
	"01111011110101",
	"01111100001110",
	"01111100100111",
	"01111101000000",
	"01111101011001",
	"01111101110010",
	"01111110001011",
	"01111110100100",
	"01111110111101",
	"01111111010110",
	"01111111101111",
	"10000000001000",
	"10000000100001",
	"10000000111010",
	"10000001010011",
	"10000001101100",
	"10000010000101",
	"10000010011110",
	"10000010110111",
	"10000011010000",
	"10000011101001",
	"10000100000010",
	"10000100011011",
	"10000100110100",
	"10000101001101",
	"10000101100110",
	"10000101111111",
	"10000110011000",
	"10000110110001",
	"10000111001010",
	"10000111100011",
	"10000111111100",
	"10001000010101",
	"10001000101110",
	"10001001000111",
	"10001001100000",
	"10001001111001",
	"10001010010010",
	"10001010101011",
	"10001011000100",
	"10001011011101",
	"10001011110110",
	"10001100001111",
	"10001100101000",
	"10001101000001",
	"10001101011010",
	"10001101110011",
	"10001110001100",
	"10001110100101",
	"10001110111110",
	"10001111010111",
	"10001111110000",
	"10010000001001",
	"10010000100010",
	"10010000111011",
	"10010001010100",
	"10010001101101",
	"10010010000110",
	"10010010011111",
	"10010010111000",
	"10010011010001",
	"10010011101010",
	"10010100000011",
	"10010100011100",
	"10010100110101",
	"10010101001110",
	"10010101100111",
	"10010110000000",
	"10010110011001",
	"10010110110010",
	"10010111001011",
	"10010111100100",
	"10010111111101",
	"10011000010110",
	"10011000101111",
	"10011001001000",
	"10011001100001",
	"10011001111010",
	"10011010010011",
	"10011010101100",
	"10011011000101",
	"10011011011110",
	"10011011110111",
	"10011100010000",
	"10011100101001",
	"10011101000010",
	"10011101011011",
	"10011101110100",
	"10011110001101",
	"10011110100110",
	"10011110111111",
	"10011111011000",
	"10011111110001",
	"10100000001010",
	"10100000100011",
	"10100000111100",
	"10100001010101",
	"10100001101110",
	"10100010000111",
	"10100010100000",
	"10100010111001",
	"10100011010010",
	"10100011101011",
	"10100100000100",
	"10100100011101",
	"10100100110110",
	"10100101001111",
	"10100101101000",
	"10100110000001",
	"10100110011010",
	"10100110110011",
	"10100111001100",
	"10100111100101",
	"10100111111110",
	"10101000010111",
	"10101000110000",
	"10101001001001",
	"10101001100010",
	"10101001111011",
	"10101010010100",
	"10101010101101",
	"10101011000110",
	"10101011011111",
	"10101011111000",
	"10101100010001",
	"10101100101010",
	"10101101000011",
	"10101101011100",
	"10101101110101",
	"10101110001110",
	"10101110100111",
	"10101111000000",
	"10101111011001",
	"10101111110010",
	"10110000001011",
	"10110000100100",
	"10110000111101",
	"10110001010110",
	"10110001101111",
	"10110010001000",
	"10110010100001",
	"10110010111010",
	"10110011010011",
	"10110011101100",
	"10110100000101",
	"10110100011110",
	"10110100110111",
	"10110101010000",
	"10110101101001",
	"10110110000010",
	"10110110011011",
	"10110110110100",
	"10110111001101",
	"10110111100110",
	"10110111111111",
	"10111000011000",
	"10111000110001",
	"10111001001010",
	"10111001100011",
	"10111001111100",
	"10111010010101",
	"10111010101110",
	"10111011000111",
	"10111011100000",
	"10111011111001",
	"10111100010010",
	"10111100101011",
	"10111101000100",
	"10111101011101",
	"10111101110110",
	"10111110001111",
	"10111110101000",
	"10111111000001",
	"10111111011010",
	"10111111110011",
	"11000000001100",
	"11000000100101",
	"11000000111110",
	"11000001010111",
	"11000001110000",
	"11000010001001",
	"11000010100010",
	"11000010111011",
	"11000011010100",
	"11000011101101",
	"11000100000110",
	"11000100011111",
	"11000100111000",
	"11000101010001",
	"11000101101010",
	"11000110000011",
	"11000110011100",
	"11000110110101",
	"11000111001110",
	"11000111100111",
	"11001000000000",
	"11001000011001",
	"11001000110010",
	"11001001001011",
	"11001001100100",
	"11001001111101",
	"11001010010110",
	"11001010101111",
	"11001011001000",
	"11001011100001",
	"11001011111010",
	"11001100010011",
	"11001100101100",
	"11001101000101",
	"11001101011110",
	"11001101110111",
	"11001110010000",
	"11001110101001",
	"11001111000010",
	"11001111011011",
	"11001111110100",
	"11010000001101",
	"11010000100110",
	"11010000111111",
	"11010001011000",
	"11010001110001",
	"11010010001010",
	"11010010100011",
	"11010010111100",
	"11010011010101",
	"11010011101110",
	"11010100000111",
	"11010100100000",
	"11010100111001",
	"11010101010010",
	"11010101101011",
	"11010110000100",
	"11010110011101",
	"11010110110110",
	"11010111001111",
	"11010111101000",
	"11011000000001",
	"11011000011010",
	"11011000110011",
	"11011001001100",
	"11011001100101",
	"11011001111110",
	"11011010010111",
	"11011010110000",
	"11011011001001",
	"11011011100010",
	"11011011111011",
	"11011100010100",
	"11011100101101",
	"11011101000110",
	"11011101011111",
	"11011101111000",
	"11011110010001",
	"11011110101010",
	"11011111000011",
	"11011111011100",
	"11011111110101",
	"11100000001110",
	"11100000100111",
	"11100001000000",
	"11100001011001",
	"11100001110010",
	"11100010001011",
	"11100010100100",
	"11100010111101",
	"11100011010110",
	"11100011101111",
	"11100100001000",
	"11100100100001",
	"11100100111010",
	"11100101010011",
	"11100101101100",
	"11100110000101",
	"11100110011110",
	"11100110110111",
	"11100111010000",
	"11100111101001",
	"11101000000010",
	"11101000011011",
	"11101000110100",
	"11101001001101",
	"11101001100110",
	"11101001111111"
);

-------------------------------------------------------------------------
-- Declare functions and procedure
-------------------------------------------------------------------------

function siga_point_to_linear (signal x : in std_logic_vector(9 downto 0);
	signal y                                : in std_logic_vector(9 downto 0)
) return std_logic_vector;
function siga_int_to_rgb (red : in integer range 0 to 31;
	green                         : in integer range 0 to 63;
	blue                          : in integer range 0 to 31
) return siga_rgb_t;

function siga_word_to_rgb (rgb : std_logic_vector(15 downto 0)
) return siga_rgb_t;

function siga_get_max (signal a : in signed;
	signal b                        : in signed
) return signed;
end package siga_utilities;

package body siga_utilities is

	function siga_point_to_linear (signal x : in std_logic_vector(9 downto 0);
		signal y                                : in std_logic_vector(9 downto 0)) return std_logic_vector is
		variable y_start_addr                   : std_logic_vector(18 downto 0);
	begin
		y_start_addr := mul_r_c_table(to_integer(unsigned(y))) & "00000";
		return std_logic_vector(unsigned(y_start_addr) + unsigned(x));
	end siga_point_to_linear;

	function siga_get_max (signal a : in signed;
		signal b                        : in signed) return signed is
	begin
		if a > b then
			return a;
		else
			return b;
		end if;
	end siga_get_max;

	function siga_int_to_rgb (red : in integer range 0 to 31;
		green                         : in integer range 0 to 63;
		blue                          : in integer range 0 to 31) return siga_rgb_t is
		variable rgb_pack             : siga_rgb_t;
	begin
		rgb_pack.r := std_logic_vector(TO_UNSIGNED(red, 5));
		rgb_pack.g := std_logic_vector(TO_UNSIGNED(green, 6));
		rgb_pack.b := std_logic_vector(TO_UNSIGNED(blue, 5));
		return rgb_pack;
	end siga_int_to_rgb;

	function siga_word_to_rgb (rgb : std_logic_vector(15 downto 0))
		return siga_rgb_t is
		variable rgb_pack : siga_rgb_t;
	begin
		rgb_pack.r := rgb(15 downto 11);
		rgb_pack.g := rgb(10 downto 5);
		rgb_pack.b := rgb(4 downto 0);
		return rgb_pack;
	end siga_word_to_rgb;

end package body siga_utilities;
